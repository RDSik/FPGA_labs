module user_not (
    input  wire a,
    output wire c
);
    assign c = ~a;

endmodule
