`timescale 1ns / 1ps  //параметры шкалы ШАГ ns / ТОЧНОСТЬ ps

module sw_led_tb ();  //название модуля тестирования

    reg [7:0] in_tb; //регистр 8 бит, выполняет роль генератора и подает значения в модуль sw_led
    wire [4:0] out_tb; //шина проводов на 5 бит, будет выполнять роль осциллографа для снятия выходных сигналов из модуля
    integer i;  //целочисленная переменная для счетчика

    sw_led DUT( //инстанцирование модуля sw_led с именем экземпляра DUT
        .in (in_tb), //подключение регистра in_tb к шине in из модуля sw_led
        .out (out_tb) //подключение шины out_tb к шине out из модуля sw_led
    );

    initial  // блок инициализации (см приложение 1)
        begin  // открытие "скобок"
            for (i = 0; i < 256; i = i + 1) begin  // открытие "скобок"
                in_tb = i; //присвоение регистру in_tb значения счетчика
                #10;
            end  // закрытие "скобок"
            $stop;
        end  // закрытие "скобок"

endmodule
