module sw_led (  //название модуля
    input  wire [7:0] in,  //входная 8-битная шина проводов
    output wire [4:0] out  //выходная 5-битная шина проводов
);

    //присвоение 4 биту шины out логической операции И между in[6] и in[7]
    assign out[4] = in[6] & in[7];
    //присвоение 3 биту шины out логической операции ИЛИ между in[5] и in[4]
    assign out[3] = in[5] | in[4];
    //присвоение 2 биту шины out логического отрицания сигнала in[3]
    assign out[2] = ~in[3];
    //присвоение 1 биту шины out логической операции И-НЕ между in[1] и in[2]
    assign out[1] = ~(in[1] & in[2]);
    //присвоение 0 биту шины out сигнала на in[0]
    assign out[0] = in[0];

endmodule  //завершение модуля
